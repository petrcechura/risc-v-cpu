

/** TODO */
interface system_bus_if(
  inout wire[15:0] IO,
  inout wire SCLK,
  inout wire ON
);
endinterface: SystemBus
